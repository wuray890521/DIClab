.SUBCKT Comparator VSS VDD  A[63] A[62] A[61] A[60] A[59] A[58] A[57] A[56] A[55] A[54] A[53] A[52] A[51] A[50] A[49] A[48] A[47] A[46] A[45] A[44] A[43] A[42] A[41] A[40] A[39] A[38] A[37] A[36] A[35] A[34] A[33] A[32] A[31] A[30] A[29] A[28] A[27] A[26] A[25] A[24] A[23] A[22] A[21] A[20] A[19] A[18] A[17] A[16] A[15] A[14] A[13] A[12] A[11] A[10] A[9] A[8] A[7] A[6] A[5] A[4] A[3] A[2] A[1] A[0] B[63] B[62] B[61] B[60] B[59] B[58] B[57] B[56] B[55] B[54] B[53] B[52] B[51] B[50] B[49] B[48] B[47] B[46] B[45] B[44] B[43] B[42] B[41] B[40] B[39] B[38] B[37] B[36] B[35] B[34] B[33] B[32] B[31] B[30] B[29] B[28] B[27] B[26] B[25] B[24] B[23] B[22] B[21] B[20] B[19] B[18] B[17] B[16] B[15] B[14] B[13] B[12] B[11] B[10] B[9] B[8] B[7] B[6] B[5] B[4] B[3] B[2] B[1] B[0] Out
XU10 VSS VDD  n1 n2 n3 n4 n5 Out NOR5xp2_ASAP7_75t_R
XU11 VSS VDD  n6 n7 n8 n9 n10 n5 NAND5xp2_ASAP7_75t_R
XU12 VSS VDD  B[4] A[4] n14 XOR2xp5_ASAP7_75t_R
XU13 VSS VDD  B[5] A[5] n13 XOR2xp5_ASAP7_75t_R
XU14 VSS VDD  B[6] A[6] n12 XOR2xp5_ASAP7_75t_R
XU15 VSS VDD  B[7] A[7] n11 XOR2xp5_ASAP7_75t_R
XU16 VSS VDD  B[3] A[3] n9 XNOR2xp5_ASAP7_75t_R
XU17 VSS VDD  B[2] A[2] n8 XNOR2xp5_ASAP7_75t_R
XU18 VSS VDD  B[1] A[1] n7 XNOR2xp5_ASAP7_75t_R
XU19 VSS VDD  B[0] A[0] n6 XNOR2xp5_ASAP7_75t_R
XU20 VSS VDD  n15 n16 n17 n18 n19 n4 NAND5xp2_ASAP7_75t_R
XU21 VSS VDD  B[14] A[14] n23 XOR2xp5_ASAP7_75t_R
XU22 VSS VDD  B[15] A[15] n22 XOR2xp5_ASAP7_75t_R
XU23 VSS VDD  B[8] A[8] n21 XOR2xp5_ASAP7_75t_R
XU24 VSS VDD  B[9] A[9] n20 XOR2xp5_ASAP7_75t_R
XU25 VSS VDD  B[13] A[13] n18 XNOR2xp5_ASAP7_75t_R
XU26 VSS VDD  B[12] A[12] n17 XNOR2xp5_ASAP7_75t_R
XU27 VSS VDD  B[11] A[11] n16 XNOR2xp5_ASAP7_75t_R
XU28 VSS VDD  B[10] A[10] n15 XNOR2xp5_ASAP7_75t_R
XU29 VSS VDD  n24 n25 n26 n27 n28 n3 NAND5xp2_ASAP7_75t_R
XU30 VSS VDD  B[20] A[20] n32 XOR2xp5_ASAP7_75t_R
XU31 VSS VDD  B[21] A[21] n31 XOR2xp5_ASAP7_75t_R
XU32 VSS VDD  B[22] A[22] n30 XOR2xp5_ASAP7_75t_R
XU33 VSS VDD  B[23] A[23] n29 XOR2xp5_ASAP7_75t_R
XU34 VSS VDD  B[19] A[19] n27 XNOR2xp5_ASAP7_75t_R
XU35 VSS VDD  B[18] A[18] n26 XNOR2xp5_ASAP7_75t_R
XU36 VSS VDD  B[17] A[17] n25 XNOR2xp5_ASAP7_75t_R
XU37 VSS VDD  B[16] A[16] n24 XNOR2xp5_ASAP7_75t_R
XU38 VSS VDD  n33 n34 n35 n36 n37 n2 NAND5xp2_ASAP7_75t_R
XU39 VSS VDD  B[36] A[36] n41 XOR2xp5_ASAP7_75t_R
XU40 VSS VDD  B[37] A[37] n40 XOR2xp5_ASAP7_75t_R
XU41 VSS VDD  B[38] A[38] n39 XOR2xp5_ASAP7_75t_R
XU42 VSS VDD  B[39] A[39] n38 XOR2xp5_ASAP7_75t_R
XU43 VSS VDD  B[35] A[35] n36 XNOR2xp5_ASAP7_75t_R
XU44 VSS VDD  B[34] A[34] n35 XNOR2xp5_ASAP7_75t_R
XU45 VSS VDD  B[33] A[33] n34 XNOR2xp5_ASAP7_75t_R
XU46 VSS VDD  B[32] A[32] n33 XNOR2xp5_ASAP7_75t_R
XU47 VSS VDD  n46 n47 n48 n49 n50 n45 NOR5xp2_ASAP7_75t_R
XU48 VSS VDD  B[24] A[24] n50 XOR2xp5_ASAP7_75t_R
XU49 VSS VDD  B[25] A[25] n49 XOR2xp5_ASAP7_75t_R
XU50 VSS VDD  B[26] A[26] n48 XOR2xp5_ASAP7_75t_R
XU51 VSS VDD  B[27] A[27] n47 XOR2xp5_ASAP7_75t_R
XU52 VSS VDD  B[31] A[31] n54 XNOR2xp5_ASAP7_75t_R
XU53 VSS VDD  B[30] A[30] n53 XNOR2xp5_ASAP7_75t_R
XU54 VSS VDD  B[29] A[29] n52 XNOR2xp5_ASAP7_75t_R
XU55 VSS VDD  B[28] A[28] n51 XNOR2xp5_ASAP7_75t_R
XU56 VSS VDD  n55 n56 n57 n58 n59 n44 NOR5xp2_ASAP7_75t_R
XU57 VSS VDD  B[56] A[56] n59 XOR2xp5_ASAP7_75t_R
XU58 VSS VDD  B[57] A[57] n58 XOR2xp5_ASAP7_75t_R
XU59 VSS VDD  B[58] A[58] n57 XOR2xp5_ASAP7_75t_R
XU60 VSS VDD  B[59] A[59] n56 XOR2xp5_ASAP7_75t_R
XU61 VSS VDD  B[63] A[63] n63 XNOR2xp5_ASAP7_75t_R
XU62 VSS VDD  B[62] A[62] n62 XNOR2xp5_ASAP7_75t_R
XU63 VSS VDD  B[61] A[61] n61 XNOR2xp5_ASAP7_75t_R
XU64 VSS VDD  B[60] A[60] n60 XNOR2xp5_ASAP7_75t_R
XU65 VSS VDD  n64 n65 n66 n67 n68 n43 NOR5xp2_ASAP7_75t_R
XU66 VSS VDD  B[48] A[48] n68 XOR2xp5_ASAP7_75t_R
XU67 VSS VDD  B[49] A[49] n67 XOR2xp5_ASAP7_75t_R
XU68 VSS VDD  B[50] A[50] n66 XOR2xp5_ASAP7_75t_R
XU69 VSS VDD  B[51] A[51] n65 XOR2xp5_ASAP7_75t_R
XU70 VSS VDD  B[55] A[55] n72 XNOR2xp5_ASAP7_75t_R
XU71 VSS VDD  B[54] A[54] n71 XNOR2xp5_ASAP7_75t_R
XU72 VSS VDD  B[53] A[53] n70 XNOR2xp5_ASAP7_75t_R
XU73 VSS VDD  B[52] A[52] n69 XNOR2xp5_ASAP7_75t_R
XU74 VSS VDD  n73 n74 n75 n76 n77 n42 NOR5xp2_ASAP7_75t_R
XU75 VSS VDD  B[40] A[40] n77 XOR2xp5_ASAP7_75t_R
XU76 VSS VDD  B[41] A[41] n76 XOR2xp5_ASAP7_75t_R
XU77 VSS VDD  B[42] A[42] n75 XOR2xp5_ASAP7_75t_R
XU78 VSS VDD  B[43] A[43] n74 XOR2xp5_ASAP7_75t_R
XU79 VSS VDD  B[47] A[47] n81 XNOR2xp5_ASAP7_75t_R
XU80 VSS VDD  B[46] A[46] n80 XNOR2xp5_ASAP7_75t_R
XU81 VSS VDD  B[45] A[45] n79 XNOR2xp5_ASAP7_75t_R
XU82 VSS VDD  B[44] A[44] n78 XNOR2xp5_ASAP7_75t_R
XU83 VSS VDD  n42 n43 n44 n45 n1 NAND4xp25_ASAP7_75t_R
XU84 VSS VDD  n60 n61 n62 n63 n55 NAND4xp25_ASAP7_75t_R
XU85 VSS VDD  n51 n52 n53 n54 n46 NAND4xp25_ASAP7_75t_R
XU86 VSS VDD  n69 n70 n71 n72 n64 NAND4xp25_ASAP7_75t_R
XU87 VSS VDD  n78 n79 n80 n81 n73 NAND4xp25_ASAP7_75t_R
XU88 VSS VDD  n11 n12 n13 n14 n10 NOR4xp25_ASAP7_75t_R
XU89 VSS VDD  n20 n21 n22 n23 n19 NOR4xp25_ASAP7_75t_R
XU90 VSS VDD  n29 n30 n31 n32 n28 NOR4xp25_ASAP7_75t_R
XU91 VSS VDD  n38 n39 n40 n41 n37 NOR4xp25_ASAP7_75t_R
Coutput1 n1 GND 3f
Coutput2 n2 GND 3f
Coutput3 n3 GND 3f
Coutput4 n4 GND 3f
Coutput5 n5 GND 3f
Coutput6 n6 GND 3f
Coutput7 n7 GND 3f
Coutput8 n8 GND 3f
Coutput9 n9 GND 3f
Coutput10 n10 GND 3f
Coutput11 n11 GND 3f
Coutput12 n12 GND 3f
Coutput13 n13 GND 3f
Coutput14 n14 GND 3f
Coutput15 n15 GND 3f
Coutput16 n16 GND 3f
Coutput17 n17 GND 3f
Coutput18 n18 GND 3f
Coutput19 n19 GND 3f
Coutput20 n20 GND 3f
Coutput21 n21 GND 3f
Coutput22 n22 GND 3f
Coutput23 n23 GND 3f
Coutput24 n24 GND 3f
Coutput25 n25 GND 3f
Coutput26 n26 GND 3f
Coutput27 n27 GND 3f
Coutput28 n28 GND 3f
Coutput29 n29 GND 3f
Coutput30 n30 GND 3f
Coutput31 n31 GND 3f
Coutput32 n32 GND 3f
Coutput33 n33 GND 3f
Coutput34 n34 GND 3f
Coutput35 n35 GND 3f
Coutput36 n36 GND 3f
Coutput37 n37 GND 3f
Coutput38 n38 GND 3f
Coutput39 n39 GND 3f
Coutput40 n40 GND 3f
Coutput41 n41 GND 3f
Coutput42 n42 GND 3f
Coutput43 n43 GND 3f
Coutput44 n44 GND 3f
Coutput45 n45 GND 3f
Coutput46 n46 GND 3f
Coutput47 n47 GND 3f
Coutput48 n48 GND 3f
Coutput49 n49 GND 3f
Coutput50 n50 GND 3f
Coutput51 n51 GND 3f
Coutput52 n52 GND 3f
Coutput53 n53 GND 3f
Coutput54 n54 GND 3f
Coutput55 n55 GND 3f
Coutput56 n56 GND 3f
Coutput57 n57 GND 3f
Coutput58 n58 GND 3f
Coutput59 n59 GND 3f
Coutput60 n60 GND 3f
Coutput61 n61 GND 3f
Coutput62 n62 GND 3f
Coutput63 n63 GND 3f
Coutput64 n64 GND 3f
Coutput65 n65 GND 3f
Coutput66 n66 GND 3f
Coutput67 n67 GND 3f
Coutput68 n68 GND 3f
Coutput69 n69 GND 3f
Coutput70 n70 GND 3f
Coutput71 n71 GND 3f
Coutput72 n72 GND 3f
Coutput73 n73 GND 3f
Coutput74 n74 GND 3f
Coutput75 n75 GND 3f
Coutput76 n76 GND 3f
Coutput77 n77 GND 3f
Coutput78 n78 GND 3f
Coutput79 n79 GND 3f
Coutput80 n80 GND 3f
Coutput81 n81 GND 3f
.ENDS


