.SUBCKT Convolution VSS VDD  IFM_0[3] IFM_0[2] IFM_0[1] IFM_0[0] IFM_1[3] IFM_1[2] IFM_1[1] IFM_1[0] IFM_2[3] IFM_2[2] IFM_2[1] IFM_2[0] IFM_3[3] IFM_3[2] IFM_3[1] IFM_3[0] INW_0[3] INW_0[2] INW_0[1] INW_0[0] INW_1[3] INW_1[2] INW_1[1] INW_1[0] INW_2[3] INW_2[2] INW_2[1] INW_2[0] INW_3[3] INW_3[2] INW_3[1] INW_3[0] Output[9] Output[8] Output[7] Output[6] Output[5] Output[4] Output[3] Output[2] Output[1] Output[0] Port10
XDP_OP_10J1_122_2300_U128 VSS VDD  DP_OP_10J1_122_2300_n203 DP_OP_10J1_122_2300_n206 DP_OP_10J1_122_2300_n227 DP_OP_10J1_122_2300_n162 DP_OP_10J1_122_2300_n163 FAx1_ASAP7_75t_R
XDP_OP_10J1_122_2300_U127 VSS VDD  DP_OP_10J1_122_2300_n230 DP_OP_10J1_122_2300_n254 DP_OP_10J1_122_2300_n251 DP_OP_10J1_122_2300_n160 DP_OP_10J1_122_2300_n161 FAx1_ASAP7_75t_R
XDP_OP_10J1_122_2300_U125 VSS VDD  DP_OP_10J1_122_2300_n165 DP_OP_10J1_122_2300_n166 DP_OP_10J1_122_2300_n157 DP_OP_10J1_122_2300_n158 DP_OP_10J1_122_2300_n159 FAx1_ASAP7_75t_R
XDP_OP_10J1_122_2300_U122 VSS VDD  DP_OP_10J1_122_2300_n175 DP_OP_10J1_122_2300_n178 DP_OP_10J1_122_2300_n181 DP_OP_10J1_122_2300_n153 DP_OP_10J1_122_2300_n154 FAx1_ASAP7_75t_R
XDP_OP_10J1_122_2300_U121 VSS VDD  DP_OP_10J1_122_2300_n199 DP_OP_10J1_122_2300_n202 DP_OP_10J1_122_2300_n205 DP_OP_10J1_122_2300_n151 DP_OP_10J1_122_2300_n152 FAx1_ASAP7_75t_R
XDP_OP_10J1_122_2300_U120 VSS VDD  DP_OP_10J1_122_2300_n223 DP_OP_10J1_122_2300_n253 DP_OP_10J1_122_2300_n226 DP_OP_10J1_122_2300_n149 DP_OP_10J1_122_2300_n150 FAx1_ASAP7_75t_R
XDP_OP_10J1_122_2300_U119 VSS VDD  DP_OP_10J1_122_2300_n229 DP_OP_10J1_122_2300_n250 DP_OP_10J1_122_2300_n247 DP_OP_10J1_122_2300_n147 DP_OP_10J1_122_2300_n148 FAx1_ASAP7_75t_R
XDP_OP_10J1_122_2300_U117 VSS VDD  DP_OP_10J1_122_2300_n162 DP_OP_10J1_122_2300_n144 DP_OP_10J1_122_2300_n160 DP_OP_10J1_122_2300_n145 DP_OP_10J1_122_2300_n146 FAx1_ASAP7_75t_R
XDP_OP_10J1_122_2300_U116 VSS VDD  DP_OP_10J1_122_2300_n152 DP_OP_10J1_122_2300_n148 DP_OP_10J1_122_2300_n154 DP_OP_10J1_122_2300_n142 DP_OP_10J1_122_2300_n143 FAx1_ASAP7_75t_R
XDP_OP_10J1_122_2300_U114 VSS VDD  DP_OP_10J1_122_2300_n158 DP_OP_10J1_122_2300_n150 DP_OP_10J1_122_2300_n139 DP_OP_10J1_122_2300_n140 DP_OP_10J1_122_2300_n141 FAx1_ASAP7_75t_R
XDP_OP_10J1_122_2300_U111 VSS VDD  DP_OP_10J1_122_2300_n177 DP_OP_10J1_122_2300_n180 DP_OP_10J1_122_2300_n195 DP_OP_10J1_122_2300_n135 DP_OP_10J1_122_2300_n136 FAx1_ASAP7_75t_R
XDP_OP_10J1_122_2300_U110 VSS VDD  DP_OP_10J1_122_2300_n198 DP_OP_10J1_122_2300_n201 DP_OP_10J1_122_2300_n204 DP_OP_10J1_122_2300_n133 DP_OP_10J1_122_2300_n134 FAx1_ASAP7_75t_R
XDP_OP_10J1_122_2300_U109 VSS VDD  DP_OP_10J1_122_2300_n219 DP_OP_10J1_122_2300_n252 DP_OP_10J1_122_2300_n222 DP_OP_10J1_122_2300_n131 DP_OP_10J1_122_2300_n132 FAx1_ASAP7_75t_R
XDP_OP_10J1_122_2300_U108 VSS VDD  DP_OP_10J1_122_2300_n225 DP_OP_10J1_122_2300_n249 DP_OP_10J1_122_2300_n228 DP_OP_10J1_122_2300_n129 DP_OP_10J1_122_2300_n130 FAx1_ASAP7_75t_R
XDP_OP_10J1_122_2300_U106 VSS VDD  DP_OP_10J1_122_2300_n243 DP_OP_10J1_122_2300_n246 DP_OP_10J1_122_2300_n126 DP_OP_10J1_122_2300_n127 DP_OP_10J1_122_2300_n128 FAx1_ASAP7_75t_R
XDP_OP_10J1_122_2300_U104 VSS VDD  DP_OP_10J1_122_2300_n147 DP_OP_10J1_122_2300_n151 DP_OP_10J1_122_2300_n123 DP_OP_10J1_122_2300_n124 DP_OP_10J1_122_2300_n125 FAx1_ASAP7_75t_R
XDP_OP_10J1_122_2300_U103 VSS VDD  DP_OP_10J1_122_2300_n132 DP_OP_10J1_122_2300_n149 DP_OP_10J1_122_2300_n130 DP_OP_10J1_122_2300_n121 DP_OP_10J1_122_2300_n122 FAx1_ASAP7_75t_R
XDP_OP_10J1_122_2300_U101 VSS VDD  DP_OP_10J1_122_2300_n136 DP_OP_10J1_122_2300_n134 DP_OP_10J1_122_2300_n118 DP_OP_10J1_122_2300_n119 DP_OP_10J1_122_2300_n120 FAx1_ASAP7_75t_R
XDP_OP_10J1_122_2300_U99 VSS VDD  DP_OP_10J1_122_2300_n142 DP_OP_10J1_122_2300_n115 DP_OP_10J1_122_2300_n125 DP_OP_10J1_122_2300_n116 DP_OP_10J1_122_2300_n117 FAx1_ASAP7_75t_R
XDP_OP_10J1_122_2300_U98 VSS VDD  DP_OP_10J1_122_2300_n120 DP_OP_10J1_122_2300_n122 DP_OP_10J1_122_2300_n140 DP_OP_10J1_122_2300_n113 DP_OP_10J1_122_2300_n114 FAx1_ASAP7_75t_R
XDP_OP_10J1_122_2300_U93 VSS VDD  DP_OP_10J1_122_2300_n176 DP_OP_10J1_122_2300_n248 DP_OP_10J1_122_2300_n194 DP_OP_10J1_122_2300_n107 DP_OP_10J1_122_2300_n108 FAx1_ASAP7_75t_R
XDP_OP_10J1_122_2300_U92 VSS VDD  DP_OP_10J1_122_2300_n197 DP_OP_10J1_122_2300_n245 DP_OP_10J1_122_2300_n200 DP_OP_10J1_122_2300_n105 DP_OP_10J1_122_2300_n106 FAx1_ASAP7_75t_R
XDP_OP_10J1_122_2300_U91 VSS VDD  DP_OP_10J1_122_2300_n218 DP_OP_10J1_122_2300_n242 DP_OP_10J1_122_2300_n221 DP_OP_10J1_122_2300_n103 DP_OP_10J1_122_2300_n104 FAx1_ASAP7_75t_R
XDP_OP_10J1_122_2300_U89 VSS VDD  DP_OP_10J1_122_2300_n137 DP_OP_10J1_122_2300_n224 DP_OP_10J1_122_2300_n100 DP_OP_10J1_122_2300_n101 DP_OP_10J1_122_2300_n102 FAx1_ASAP7_75t_R
XDP_OP_10J1_122_2300_U87 VSS VDD  DP_OP_10J1_122_2300_n129 DP_OP_10J1_122_2300_n133 DP_OP_10J1_122_2300_n97 DP_OP_10J1_122_2300_n98 DP_OP_10J1_122_2300_n99 FAx1_ASAP7_75t_R
XDP_OP_10J1_122_2300_U86 VSS VDD  DP_OP_10J1_122_2300_n104 DP_OP_10J1_122_2300_n131 DP_OP_10J1_122_2300_n106 DP_OP_10J1_122_2300_n95 DP_OP_10J1_122_2300_n96 FAx1_ASAP7_75t_R
XDP_OP_10J1_122_2300_U84 VSS VDD  DP_OP_10J1_122_2300_n127 DP_OP_10J1_122_2300_n108 DP_OP_10J1_122_2300_n92 DP_OP_10J1_122_2300_n93 DP_OP_10J1_122_2300_n94 FAx1_ASAP7_75t_R
XDP_OP_10J1_122_2300_U82 VSS VDD  DP_OP_10J1_122_2300_n89 DP_OP_10J1_122_2300_n121 DP_OP_10J1_122_2300_n99 DP_OP_10J1_122_2300_n90 DP_OP_10J1_122_2300_n91 FAx1_ASAP7_75t_R
XDP_OP_10J1_122_2300_U80 VSS VDD  DP_OP_10J1_122_2300_n96 DP_OP_10J1_122_2300_n119 DP_OP_10J1_122_2300_n86 DP_OP_10J1_122_2300_n87 DP_OP_10J1_122_2300_n88 FAx1_ASAP7_75t_R
XDP_OP_10J1_122_2300_U78 VSS VDD  DP_OP_10J1_122_2300_n91 DP_OP_10J1_122_2300_n83 DP_OP_10J1_122_2300_n113 DP_OP_10J1_122_2300_n84 DP_OP_10J1_122_2300_n85 FAx1_ASAP7_75t_R
XDP_OP_10J1_122_2300_U74 VSS VDD  DP_OP_10J1_122_2300_n172 DP_OP_10J1_122_2300_n241 DP_OP_10J1_122_2300_n193 DP_OP_10J1_122_2300_n78 DP_OP_10J1_122_2300_n79 FAx1_ASAP7_75t_R
XDP_OP_10J1_122_2300_U73 VSS VDD  DP_OP_10J1_122_2300_n196 DP_OP_10J1_122_2300_n220 DP_OP_10J1_122_2300_n217 DP_OP_10J1_122_2300_n76 DP_OP_10J1_122_2300_n77 FAx1_ASAP7_75t_R
XDP_OP_10J1_122_2300_U71 VSS VDD  DP_OP_10J1_122_2300_n107 DP_OP_10J1_122_2300_n73 DP_OP_10J1_122_2300_n105 DP_OP_10J1_122_2300_n74 DP_OP_10J1_122_2300_n75 FAx1_ASAP7_75t_R
XDP_OP_10J1_122_2300_U69 VSS VDD  DP_OP_10J1_122_2300_n70 DP_OP_10J1_122_2300_n103 DP_OP_10J1_122_2300_n77 DP_OP_10J1_122_2300_n71 DP_OP_10J1_122_2300_n72 FAx1_ASAP7_75t_R
XDP_OP_10J1_122_2300_U67 VSS VDD  DP_OP_10J1_122_2300_n101 DP_OP_10J1_122_2300_n79 DP_OP_10J1_122_2300_n67 DP_OP_10J1_122_2300_n68 DP_OP_10J1_122_2300_n69 FAx1_ASAP7_75t_R
XDP_OP_10J1_122_2300_U66 VSS VDD  DP_OP_10J1_122_2300_n75 DP_OP_10J1_122_2300_n95 DP_OP_10J1_122_2300_n93 DP_OP_10J1_122_2300_n65 DP_OP_10J1_122_2300_n66 FAx1_ASAP7_75t_R
XDP_OP_10J1_122_2300_U64 VSS VDD  DP_OP_10J1_122_2300_n69 DP_OP_10J1_122_2300_n72 DP_OP_10J1_122_2300_n62 DP_OP_10J1_122_2300_n63 DP_OP_10J1_122_2300_n64 FAx1_ASAP7_75t_R
XDP_OP_10J1_122_2300_U62 VSS VDD  DP_OP_10J1_122_2300_n87 DP_OP_10J1_122_2300_n66 DP_OP_10J1_122_2300_n59 DP_OP_10J1_122_2300_n60 DP_OP_10J1_122_2300_n61 FAx1_ASAP7_75t_R
XDP_OP_10J1_122_2300_U58 VSS VDD  DP_OP_10J1_122_2300_n192 DP_OP_10J1_122_2300_n216 DP_OP_10J1_122_2300_n80 DP_OP_10J1_122_2300_n54 DP_OP_10J1_122_2300_n55 FAx1_ASAP7_75t_R
XDP_OP_10J1_122_2300_U56 VSS VDD  DP_OP_10J1_122_2300_n76 DP_OP_10J1_122_2300_n78 DP_OP_10J1_122_2300_n51 DP_OP_10J1_122_2300_n52 DP_OP_10J1_122_2300_n53 FAx1_ASAP7_75t_R
XDP_OP_10J1_122_2300_U54 VSS VDD  DP_OP_10J1_122_2300_n48 DP_OP_10J1_122_2300_n74 DP_OP_10J1_122_2300_n71 DP_OP_10J1_122_2300_n49 DP_OP_10J1_122_2300_n50 FAx1_ASAP7_75t_R
XDP_OP_10J1_122_2300_U52 VSS VDD  DP_OP_10J1_122_2300_n68 DP_OP_10J1_122_2300_n53 DP_OP_10J1_122_2300_n45 DP_OP_10J1_122_2300_n46 DP_OP_10J1_122_2300_n47 FAx1_ASAP7_75t_R
XDP_OP_10J1_122_2300_U51 VSS VDD  DP_OP_10J1_122_2300_n63 DP_OP_10J1_122_2300_n50 DP_OP_10J1_122_2300_n47 DP_OP_10J1_122_2300_n43 DP_OP_10J1_122_2300_n44 FAx1_ASAP7_75t_R
XDP_OP_10J1_122_2300_U49 VSS VDD  DP_OP_10J1_122_2300_n40 DP_OP_10J1_122_2300_n56 DP_OP_10J1_122_2300_n52 DP_OP_10J1_122_2300_n41 DP_OP_10J1_122_2300_n42 FAx1_ASAP7_75t_R
XDP_OP_10J1_122_2300_U48 VSS VDD  DP_OP_10J1_122_2300_n42 DP_OP_10J1_122_2300_n49 DP_OP_10J1_122_2300_n46 DP_OP_10J1_122_2300_n38 DP_OP_10J1_122_2300_n39 FAx1_ASAP7_75t_R
XU1 VSS VDD  DP_OP_10J1_122_2300_n84 DP_OP_10J1_122_2300_n59 INVxp33_ASAP7_75t_R
XU2 VSS VDD  DP_OP_10J1_122_2300_n102 DP_OP_10J1_122_2300_n89 INVxp67_ASAP7_75t_R
XU3 VSS VDD  INW_0[1] n26 INVxp67_ASAP7_75t_R
XU4 VSS VDD  DP_OP_10J1_122_2300_n61 n51 INVx1_ASAP7_75t_R
XU5 VSS VDD  DP_OP_10J1_122_2300_n85 n1 HB1xp67_ASAP7_75t_R
XU6 VSS VDD  INW_2[3] IFM_2[3] n60 NAND2xp33_ASAP7_75t_R
XU7 VSS VDD  IFM_3[3] INW_3[3] n61 NAND2xp33_ASAP7_75t_R
XU8 VSS VDD  IFM_0[1] n23 INVxp33_ASAP7_75t_R
XU9 VSS VDD  INW_0[0] n38 INVxp33_ASAP7_75t_R
XU10 VSS VDD  IFM_3[0] n35 INVxp33_ASAP7_75t_R
XU11 VSS VDD  INW_3[0] n36 INVxp33_ASAP7_75t_R
XU12 VSS VDD  IFM_0[0] n37 INVxp33_ASAP7_75t_R
XU13 VSS VDD  INW_3[1] IFM_3[2] n5 NAND2xp33_ASAP7_75t_R
XU14 VSS VDD  INW_3[0] IFM_3[3] n6 NAND2xp33_ASAP7_75t_R
XU15 VSS VDD  DP_OP_10J1_122_2300_n153 DP_OP_10J1_122_2300_n126 INVxp33_ASAP7_75t_R
XU16 VSS VDD  DP_OP_10J1_122_2300_n65 DP_OP_10J1_122_2300_n45 INVxp33_ASAP7_75t_R
XU17 VSS VDD  DP_OP_10J1_122_2300_n55 DP_OP_10J1_122_2300_n48 INVxp33_ASAP7_75t_R
XU18 VSS VDD  INW_1[0] IFM_1[0] n40 NAND2xp33_ASAP7_75t_R
XU19 VSS VDD  DP_OP_10J1_122_2300_n88 n50 INVxp33_ASAP7_75t_R
XU20 VSS VDD  DP_OP_10J1_122_2300_n90 DP_OP_10J1_122_2300_n62 INVxp33_ASAP7_75t_R
XU21 VSS VDD  DP_OP_10J1_122_2300_n54 DP_OP_10J1_122_2300_n40 INVxp33_ASAP7_75t_R
XU22 VSS VDD  INW_2[3] n29 INVxp33_ASAP7_75t_R
XU23 VSS VDD  INW_3[3] n11 INVxp33_ASAP7_75t_R
XU24 VSS VDD  INW_2[2] n32 INVxp33_ASAP7_75t_R
XU25 VSS VDD  IFM_0[2] n22 INVxp33_ASAP7_75t_R
XU26 VSS VDD  INW_1[2] n18 INVxp33_ASAP7_75t_R
XU27 VSS VDD  IFM_1[2] n14 INVxp33_ASAP7_75t_R
XU28 VSS VDD  INW_0[2] n25 INVxp33_ASAP7_75t_R
XU29 VSS VDD  IFM_3[2] n9 INVxp33_ASAP7_75t_R
XU30 VSS VDD  IFM_2[2] n28 INVxp33_ASAP7_75t_R
XU31 VSS VDD  IFM_2[3] n27 INVxp33_ASAP7_75t_R
XU32 VSS VDD  DP_OP_10J1_122_2300_n135 DP_OP_10J1_122_2300_n100 INVxp33_ASAP7_75t_R
XU33 VSS VDD  n3 n2 n4 NAND2xp33_ASAP7_75t_R
XU34 VSS VDD  IFM_3[3] INW_3[1] n3 NAND2xp33_ASAP7_75t_R
XU35 VSS VDD  IFM_0[3] n21 INVxp33_ASAP7_75t_R
XU36 VSS VDD  INW_0[3] n24 INVxp33_ASAP7_75t_R
XU37 VSS VDD  INW_1[3] n17 INVxp33_ASAP7_75t_R
XU38 VSS VDD  IFM_1[3] n13 INVxp33_ASAP7_75t_R
XU39 VSS VDD  IFM_2[1] n30 INVxp33_ASAP7_75t_R
XU40 VSS VDD  IFM_3[0] INW_3[1] n8 NAND2xp33_ASAP7_75t_R
XU41 VSS VDD  INW_3[0] IFM_3[1] n7 NAND2xp33_ASAP7_75t_R
XU42 VSS VDD  INW_2[0] n31 INVxp33_ASAP7_75t_R
XU43 VSS VDD  INW_2[3] IFM_2[2] n62 NAND2xp33_ASAP7_75t_R
XU44 VSS VDD  IFM_3[3] INW_3[2] n63 NAND2xp33_ASAP7_75t_R
XU45 VSS VDD  n41 n42 INVxp33_ASAP7_75t_R
XU46 VSS VDD  DP_OP_10J1_122_2300_n146 DP_OP_10J1_122_2300_n139 INVxp33_ASAP7_75t_R
XU47 VSS VDD  DP_OP_10J1_122_2300_n128 DP_OP_10J1_122_2300_n115 INVxp33_ASAP7_75t_R
XU48 VSS VDD  n54 n53 INVxp33_ASAP7_75t_R
XU49 VSS VDD  n56 n55 INVxp33_ASAP7_75t_R
XU50 VSS VDD  DP_OP_10J1_122_2300_n38 n59 INVxp33_ASAP7_75t_R
XU51 VSS VDD  IFM_3[2] INW_3[2] n2 NAND2xp33_ASAP7_75t_R
XU52 VSS VDD  IFM_3[1] n10 INVxp33_ASAP7_75t_R
XU53 VSS VDD  INW_3[2] n12 INVxp33_ASAP7_75t_R
XU54 VSS VDD  n4 DP_OP_10J1_122_2300_n73 DP_OP_10J1_122_2300_n97 NAND2xp33_ASAP7_75t_R
XU55 VSS VDD  DP_OP_10J1_122_2300_n124 DP_OP_10J1_122_2300_n92 INVxp33_ASAP7_75t_R
XU56 VSS VDD  DP_OP_10J1_122_2300_n145 DP_OP_10J1_122_2300_n118 INVxp33_ASAP7_75t_R
XU57 VSS VDD  DP_OP_10J1_122_2300_n98 DP_OP_10J1_122_2300_n67 INVxp33_ASAP7_75t_R
XU58 VSS VDD  INW_2[0] IFM_2[0] n39 NAND2xp33_ASAP7_75t_R
XU59 VSS VDD  DP_OP_10J1_122_2300_n163 DP_OP_10J1_122_2300_n157 INVxp33_ASAP7_75t_R
XU60 VSS VDD  DP_OP_10J1_122_2300_n94 DP_OP_10J1_122_2300_n83 INVxp33_ASAP7_75t_R
XU61 VSS VDD  n47 n46 INVxp33_ASAP7_75t_R
XU62 VSS VDD  DP_OP_10J1_122_2300_n116 DP_OP_10J1_122_2300_n86 INVx1_ASAP7_75t_R
XU63 VSS VDD  IFM_3[3] INW_3[1] IFM_3[2] INW_3[2] DP_OP_10J1_122_2300_n73 NAND4xp25_ASAP7_75t_R
XU64 VSS VDD  IFM_2[0] n34 INVx1_ASAP7_75t_R
XU65 VSS VDD  n34 n29 DP_OP_10J1_122_2300_n252 NOR2xp33_ASAP7_75t_R
XU66 VSS VDD  n38 n21 DP_OP_10J1_122_2300_n219 NOR2xp33_ASAP7_75t_R
XU67 VSS VDD  n6 n5 A0  DP_OP_10J1_122_2300_n123 HAxp5_ASAP7_75t_R
XU68 VSS VDD  INW_3[0] IFM_3[3] INW_3[1] IFM_3[2] DP_OP_10J1_122_2300_n137 AND4x1_ASAP7_75t_R
XU69 VSS VDD  INW_3[0] IFM_3[0] INW_3[1] IFM_3[1] DP_OP_10J1_122_2300_n144 NAND4xp25_ASAP7_75t_R
XU70 VSS VDD  n8 n7 DP_OP_10J1_122_2300_n165 XOR2xp5_ASAP7_75t_R
XU71 VSS VDD  INW_1[0] n16 INVx1_ASAP7_75t_R
XU72 VSS VDD  IFM_1[0] n20 INVx1_ASAP7_75t_R
XU73 VSS VDD  n16 n20 n31 n34 DP_OP_10J1_122_2300_n166 NOR4xp25_ASAP7_75t_R
XU74 VSS VDD  n9 n11 DP_OP_10J1_122_2300_n172 NOR2xp33_ASAP7_75t_R
XU75 VSS VDD  n36 n9 DP_OP_10J1_122_2300_n175 NOR2xp33_ASAP7_75t_R
XU76 VSS VDD  n10 n11 DP_OP_10J1_122_2300_n176 NOR2xp33_ASAP7_75t_R
XU77 VSS VDD  n10 n12 DP_OP_10J1_122_2300_n177 NOR2xp33_ASAP7_75t_R
XU78 VSS VDD  INW_3[1] IFM_3[1] DP_OP_10J1_122_2300_n178 AND2x2_ASAP7_75t_R
XU79 VSS VDD  n35 n11 DP_OP_10J1_122_2300_n180 NOR2xp33_ASAP7_75t_R
XU80 VSS VDD  n35 n12 DP_OP_10J1_122_2300_n181 NOR2xp33_ASAP7_75t_R
XU81 VSS VDD  n17 n13 DP_OP_10J1_122_2300_n192 NOR2xp33_ASAP7_75t_R
XU82 VSS VDD  n13 n18 DP_OP_10J1_122_2300_n193 NOR2xp33_ASAP7_75t_R
XU83 VSS VDD  INW_1[1] n19 INVx1_ASAP7_75t_R
XU84 VSS VDD  n13 n19 DP_OP_10J1_122_2300_n194 NOR2xp33_ASAP7_75t_R
XU85 VSS VDD  n16 n13 DP_OP_10J1_122_2300_n195 NOR2xp33_ASAP7_75t_R
XU86 VSS VDD  n17 n14 DP_OP_10J1_122_2300_n196 NOR2xp33_ASAP7_75t_R
XU87 VSS VDD  n18 n14 DP_OP_10J1_122_2300_n197 NOR2xp33_ASAP7_75t_R
XU88 VSS VDD  n19 n14 DP_OP_10J1_122_2300_n198 NOR2xp33_ASAP7_75t_R
XU89 VSS VDD  n16 n14 DP_OP_10J1_122_2300_n199 NOR2xp33_ASAP7_75t_R
XU90 VSS VDD  IFM_1[1] n15 INVx1_ASAP7_75t_R
XU91 VSS VDD  n17 n15 DP_OP_10J1_122_2300_n200 NOR2xp33_ASAP7_75t_R
XU92 VSS VDD  n18 n15 DP_OP_10J1_122_2300_n201 NOR2xp33_ASAP7_75t_R
XU93 VSS VDD  n19 n15 DP_OP_10J1_122_2300_n202 NOR2xp33_ASAP7_75t_R
XU94 VSS VDD  n16 n15 DP_OP_10J1_122_2300_n203 NOR2xp33_ASAP7_75t_R
XU95 VSS VDD  n20 n17 DP_OP_10J1_122_2300_n204 NOR2xp33_ASAP7_75t_R
XU96 VSS VDD  n20 n18 DP_OP_10J1_122_2300_n205 NOR2xp33_ASAP7_75t_R
XU97 VSS VDD  n20 n19 DP_OP_10J1_122_2300_n206 NOR2xp33_ASAP7_75t_R
XU98 VSS VDD  n24 n21 DP_OP_10J1_122_2300_n216 NOR2xp33_ASAP7_75t_R
XU99 VSS VDD  n21 n25 DP_OP_10J1_122_2300_n217 NOR2xp33_ASAP7_75t_R
XU100 VSS VDD  n21 n26 DP_OP_10J1_122_2300_n218 NOR2xp33_ASAP7_75t_R
XU101 VSS VDD  n24 n22 DP_OP_10J1_122_2300_n220 NOR2xp33_ASAP7_75t_R
XU102 VSS VDD  n25 n22 DP_OP_10J1_122_2300_n221 NOR2xp33_ASAP7_75t_R
XU103 VSS VDD  n26 n22 DP_OP_10J1_122_2300_n222 NOR2xp33_ASAP7_75t_R
XU104 VSS VDD  n38 n22 DP_OP_10J1_122_2300_n223 NOR2xp33_ASAP7_75t_R
XU105 VSS VDD  n24 n23 DP_OP_10J1_122_2300_n224 NOR2xp33_ASAP7_75t_R
XU106 VSS VDD  n25 n23 DP_OP_10J1_122_2300_n225 NOR2xp33_ASAP7_75t_R
XU107 VSS VDD  n26 n23 DP_OP_10J1_122_2300_n226 NOR2xp33_ASAP7_75t_R
XU108 VSS VDD  n38 n23 DP_OP_10J1_122_2300_n227 NOR2xp33_ASAP7_75t_R
XU109 VSS VDD  n37 n24 DP_OP_10J1_122_2300_n228 NOR2xp33_ASAP7_75t_R
XU110 VSS VDD  n37 n25 DP_OP_10J1_122_2300_n229 NOR2xp33_ASAP7_75t_R
XU111 VSS VDD  n37 n26 DP_OP_10J1_122_2300_n230 NOR2xp33_ASAP7_75t_R
XU112 VSS VDD  n27 n32 DP_OP_10J1_122_2300_n241 NOR2xp33_ASAP7_75t_R
XU113 VSS VDD  INW_2[1] n33 INVx1_ASAP7_75t_R
XU114 VSS VDD  n27 n33 DP_OP_10J1_122_2300_n242 NOR2xp33_ASAP7_75t_R
XU115 VSS VDD  n31 n27 DP_OP_10J1_122_2300_n243 NOR2xp33_ASAP7_75t_R
XU116 VSS VDD  n28 n32 DP_OP_10J1_122_2300_n245 NOR2xp33_ASAP7_75t_R
XU117 VSS VDD  n28 n33 DP_OP_10J1_122_2300_n246 NOR2xp33_ASAP7_75t_R
XU118 VSS VDD  n31 n28 DP_OP_10J1_122_2300_n247 NOR2xp33_ASAP7_75t_R
XU119 VSS VDD  n29 n30 DP_OP_10J1_122_2300_n248 NOR2xp33_ASAP7_75t_R
XU120 VSS VDD  n32 n30 DP_OP_10J1_122_2300_n249 NOR2xp33_ASAP7_75t_R
XU121 VSS VDD  n33 n30 DP_OP_10J1_122_2300_n250 NOR2xp33_ASAP7_75t_R
XU122 VSS VDD  n31 n30 DP_OP_10J1_122_2300_n251 NOR2xp33_ASAP7_75t_R
XU123 VSS VDD  n34 n32 DP_OP_10J1_122_2300_n253 NOR2xp33_ASAP7_75t_R
XU124 VSS VDD  n34 n33 DP_OP_10J1_122_2300_n254 NOR2xp33_ASAP7_75t_R
XU125 VSS VDD  n36 n35 n44 NOR2xp33_ASAP7_75t_R
XU126 VSS VDD  n38 n37 n43 NOR2xp33_ASAP7_75t_R
XU127 VSS VDD  n40 n39 A1  n41 HAxp5_ASAP7_75t_R
XU128 VSS VDD  n44 n43 n41 A2  Output[0] FAx1_ASAP7_75t_R
XU129 VSS VDD  n44 n43 n42 n45 MAJIxp5_ASAP7_75t_R
XU130 VSS VDD  DP_OP_10J1_122_2300_n159 DP_OP_10J1_122_2300_n161 n45 A3  Output[1] FAx1_ASAP7_75t_R
XU131 VSS VDD  DP_OP_10J1_122_2300_n159 DP_OP_10J1_122_2300_n161 n45 n47 MAJIxp5_ASAP7_75t_R
XU132 VSS VDD  DP_OP_10J1_122_2300_n141 n46 DP_OP_10J1_122_2300_n143 A4  Output[2] FAx1_ASAP7_75t_R
XU133 VSS VDD  DP_OP_10J1_122_2300_n141 DP_OP_10J1_122_2300_n143 n47 n48 MAJIxp5_ASAP7_75t_R
XU134 VSS VDD  DP_OP_10J1_122_2300_n114 DP_OP_10J1_122_2300_n117 n48 A5  Output[3] FAx1_ASAP7_75t_R
XU135 VSS VDD  DP_OP_10J1_122_2300_n114 DP_OP_10J1_122_2300_n117 n48 n49 MAJIxp5_ASAP7_75t_R
XU136 VSS VDD  n1 DP_OP_10J1_122_2300_n88 n49 A6  Output[4] FAx1_ASAP7_75t_R
XU137 VSS VDD  n1 n50 n49 n52 MAJIxp5_ASAP7_75t_R
XU138 VSS VDD  DP_OP_10J1_122_2300_n64 n52 n51 A7  Output[5] FAx1_ASAP7_75t_R
XU139 VSS VDD  DP_OP_10J1_122_2300_n64 n52 n51 n54 MAJIxp5_ASAP7_75t_R
XU140 VSS VDD  DP_OP_10J1_122_2300_n60 n53 DP_OP_10J1_122_2300_n44 A8  Output[6] FAx1_ASAP7_75t_R
XU141 VSS VDD  DP_OP_10J1_122_2300_n60 DP_OP_10J1_122_2300_n44 n54 n56 MAJx2_ASAP7_75t_R
XU142 VSS VDD  DP_OP_10J1_122_2300_n39 n55 DP_OP_10J1_122_2300_n43 A9  Output[7] FAx1_ASAP7_75t_R
XU143 VSS VDD  DP_OP_10J1_122_2300_n39 DP_OP_10J1_122_2300_n43 n56 n58 MAJIxp5_ASAP7_75t_R
XU144 VSS VDD  n58 n57 INVx1_ASAP7_75t_R
XU145 VSS VDD  DP_OP_10J1_122_2300_n38 n57 DP_OP_10J1_122_2300_n41 A10  Output[8] FAx1_ASAP7_75t_R
XU146 VSS VDD  DP_OP_10J1_122_2300_n41 n59 n58 Output[9] MAJIxp5_ASAP7_75t_R
XU147 VSS VDD  n61 n60 A11  DP_OP_10J1_122_2300_n51 HAxp5_ASAP7_75t_R
XU148 VSS VDD  IFM_3[3] INW_3[3] INW_2[3] IFM_2[3] DP_OP_10J1_122_2300_n56 AND4x1_ASAP7_75t_R
XU149 VSS VDD  n63 n62 A12  DP_OP_10J1_122_2300_n70 HAxp5_ASAP7_75t_R
XU150 VSS VDD  IFM_3[3] INW_2[3] INW_3[2] IFM_2[2] DP_OP_10J1_122_2300_n80 AND4x1_ASAP7_75t_R
.ENDS


